module FSM()