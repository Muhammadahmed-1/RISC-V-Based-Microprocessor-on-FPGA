module topmodule()